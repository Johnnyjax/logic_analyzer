-- Listing 13.1
-- ROM with synchonous read (inferring Block RAM)
-- character ROM
--   - 8-by-16 (8-by-2^4) font
--   - 128 (2^7) characters
--   - ROM size: 512-by-8 (2^11-by-8) bits
--               16K bits: 1 BRAM

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity font_rom is
   port(
      clk: in std_logic;
      addr: in std_logic_vector(6 downto 0);
      data: out std_logic_vector(7 downto 0)
   );
end font_rom;

architecture arch of font_rom is
   constant ADDR_WIDTH: integer:=7;
   constant DATA_WIDTH: integer:=8;
   signal data_reg: std_logic_vector(DATA_WIDTH-1 downto 0);
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant ROM: rom_type:=(   -- 2^11-by-8
    
	"00000000", 
   "00000000", 
   "00000000",
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
	"00000000", 
   "00000000", 
   "00000000",
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "11111111", 
   "11111111", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
	
	"00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
	"00011111",
	"00011111",
	"00011000", 
	"00011000",
	"00011000", 
	"00011000",
	"00011000",
	"00011000",
	"00011000",
   "00011000", 
	"00011000",
	"00011000",
	"00011000",
   "00011000", 
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000", 
	"00011000",
	"00011000",
	"00011000",
	"11111000",
	"11111000",
   "00000000", 
	"00000000",
	"00000000",
	"00000000", 
	
	"00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
	"11111000",
	"11111000",
	"00011000", 
	"00011000",
	"00011000",
	"00011000",
	"00011000",
   "00011000", 
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000", 
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000",
	"00011000", 
	"00011000",
	"00011111",
	"00011111",
   "00000000", 
	"00000000",
	"00000000",
	"00000000",
	
	"00000000", 
   "00000000", 
   "00000000",
   "00000000", 
   "11111111", 
   "11111111", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
	"00000000", 
   "00000000", 
   "00000000",
   "00000000", 
   "00000000", 
	"00000000", 
   "00000000", 
   "00000000",
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000", 
   "00000000"
	);
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (clk'event and clk = '1') then
        data_reg <= ROM(to_integer(unsigned(addr)));
      end if;
   end process;
   data <= data_reg;
end arch;

